typedef enum { UVM_PASSIVE,UVM_ACTIVE} is_active_passive ;
